library verilog;
use verilog.vl_types.all;
entity experiment4a_v_unit is
end experiment4a_v_unit;
