library verilog;
use verilog.vl_types.all;
entity tb_experiment4a_v_unit is
end tb_experiment4a_v_unit;
