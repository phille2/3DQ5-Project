library verilog;
use verilog.vl_types.all;
entity SRAM_BIST_v_unit is
end SRAM_BIST_v_unit;
